module calculadora(
  input   [7:0] entrada_A,
  input   [7:0] entrada_B,
  input   [2:0] codigo,
  output  [7:0] saida
);

// insira seu código aqui

assign saida =   (codigo == 3'b000) ? 8'b00000000 :       // zerar
                 (codigo == 3'b001) ? entrada_A    :      // mostrar A
                 (codigo == 3'b010) ? entrada_B    :      // mostrar B
                 (codigo == 3'b011) ? entrada_A + entrada_B : // somar
                 (codigo == 3'b100) ? entrada_A - entrada_B : // subtrair
                 8'b00000000; // padrão para códigos inválidos


endmodule
